// <h1>An in-class exercise on timers</h1>
module micro(
    input clk,
    output [7:0] pc,
    output [7:0] w
);

endmodule
