// <h1><code>in-class.v</code> - skeleton code for in-class exercises</h1>
module in_class(
    input a,
    input b,
    output y
);
    assign y = a & b;

endmodule
