`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
module lab5dpath(x1,x2,x3,y,clk);
input clk;
input [9:0] x1,x2,x3;
output [9:0] y;


 
endmodule

