// # `in-class.v` - skeleton code for in-class exercises
module in_class(
    input a,
    input b,
    output y
);
    assign y = a & b;

endmodule
