// <h1>An in-class exercise on timers</h1>
module timer(
    input clk,
    input [15:0] din,
    input ld,
    input cnt_end,
	input aclr,
    output [15:0] dout
);

endmodule
