// # `in-class.v` - skeleton code for in-class exercises
module in_class(
    input logic a,
    input logic b,
    output logic y
);
    assign y = a & b;

endmodule
